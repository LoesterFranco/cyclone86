/* ---------------------------------------------------------------------
 * Центральный исполнительно-декодирующий модуль
 * Принимает на вход данные с загружаемого кодового буфера,
 * интерпретирует префиксы, опкоды, modrm, immediate и вычисляет
 * итоговые результаты, а также устанавливает необходимые запросы к
 * памяти или данным
 * ------------------------------------------------------------------ */

module decoder
(
    // Данные для анализа и декодера
    input   wire [127:0]    i_codebuf,  // Исходный даннее
    input   wire [  1:0]    align       // При невыровненных

    // Входящий регистровый файл
);

// Шаг 0 .Выравнивание кода, если данные не были выровнены ранее (0-3 байта)
wire [127:0] a_codebuf = align[0] ? i_codebuf[127: 8] : i_codebuf;
wire [127:0] b_codebuf = align[1] ? a_codebuf[127:16] : a_codebuf;

// Шаг 1. Декодирование до 3-х префиксов
`include "prefix.v"

// Шаг 2. Удаление префиксов из кодового буфера
wire [127:0] c_codebuf = p_size[0] ? b_codebuf[127: 8] : b_codebuf;
wire [127:0]   codebuf = p_size[1] ? c_codebuf[127:16] : c_codebuf;


// Декодирование опкода и наличия байта modrm, зависит от префиксов
// Декодирование modrm
// Декодирование immediate
// Вычисление результата (в том числе возможен вход из общей памяти)
// Выдача запросов на память, если есть, ea, и прочего, что нужно сделать
// -- на следующих тактах, т.е. досбор данных

endmodule
